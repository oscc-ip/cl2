
module cl2_tcm();

endmodule