`ifndef CL2_ARCH_DESC_SVH
`define CL2_ARCH_DESC_SVH

`define CL2_XLEN          32
`define CL2_REGFILE_NUM   32 // NOTE: just for I extension
`define CL2_REGFILE_WIDTH $clog2(`CL2_REGFILE_NUM)

`endif 