`include "cl2_arch_desc.svh"

module cl2_idu_i_extn(

);


endmodule