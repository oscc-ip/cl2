
module cl2_pl_ifu ();
endmodule
