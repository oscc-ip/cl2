module cl2_pl_ifu_bpu ();
endmodule
