`ifndef CL2_ARCH_DESC_SVH
`define CL2_ARCH_DESC_SVH

`define CL2_REGFILE_WIDTH 5
`define CL2_XLEN          32
`define CL2_REGFILE_NUM   32

`endif 