module cl2_pl_ifu_tinyidu #() ();

endmodule
