module cl2_rcu ();
endmodule
